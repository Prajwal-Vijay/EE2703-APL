R1   2 GND 1
V1   1 GND dc 4
V2   1 2 dc 3
.circuit
R1 n1 GND 1
R2 n2 n1 2
R3 n2 n1 3
V1 n3 n2 dc 1
.end